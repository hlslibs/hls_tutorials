/home/dgb/sb/sif/subprojs/sif_toolkits/any/Isrc/training/WalkThroughs/ImageProcessing/SlidingWindow/ram_1k_16_sp.vhd